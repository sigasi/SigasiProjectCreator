package testpackage is
	
end package testpackage;

package body testpackage is
	
end package body testpackage;
