package foo is
	
end package foo;

package body foo is
	
end package body foo;
